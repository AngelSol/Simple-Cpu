library verilog;
use verilog.vl_types.all;
entity outreg_vlg_vec_tst is
end outreg_vlg_vec_tst;
